module datapath_proc (clk, resetn);

	input clk, resetn;
	
	wire [15:0] NPC_IF, NPC_ID, NPC_RD, NPC_EX, NPC_MEM, NPC_WB;
	wire [15:0] PC_IF, PC_ID, PC_RD, PC_EX, PC_MEM, PC_WB;
	wire [15:0] IR_IF, IR_ID;
	
	//ID_RD
	wire [2:0] REG1ADD_ID, REG2ADD_ID, REG3ADD_ID, REG1ADD_RD, REG2ADD_RD, REG3ADD_RD;
	wire REGWRITE_ID,MEMTOREG_ID,MEMREAD_ID,MEMWRITE_ID,BRANCH_ID,REGDEST_ID, 
			REGWRITE_RD,MEMTOREG_RD,MEMREAD_RD,MEMWRITE_RD,BRANCH_RD,REGDEST_RD;
	wire [1:0] ALUSRC_ID, ALUSRC_RD;
	wire [3:0] ALUOP_ID;
	wire [5:0] IMM6_ID, IMM6_RD, IMM6_EX;
	
	//RD_EX
	wire [15:0] REG1DATA_RD, REG2DATA_RD, REG1DATA_EX, REG2DATA_EX;
	wire [2:0] REGDST_RD, REGDST_EX;
	wire REGWRITE_EX,MEMTOREG_EX,MEMREAD_EX,MEMWRITE_EX,BRANCH_EX;
	wire [1:0] ALUSRC_EX;
	wire [3:0] ALUOP_RD, ALUOP_EX;
	
	//EX_MEM
	wire ALU_Z_EX, ALU_Z_MEM, ALU_C_EX, ALU_C_MEM;
	wire [15:0] ALU_RESULT_EX, ALU_RESULT_MEM, REG2DATA_MEM;
	wire [2:0] REGDST_MEM;
	wire REGWRITE_MEM, MEMTOREG_MEM, MEMREAD_MEM, MEMWRITE_MEM, BRANCH_MEM;	
			
	//MEM_WB
	wire [15:0] MEMRD_DATA_MEM, MEMRD_DATA_WB, ALU_RESULT_WB;
	wire [2:0] REGDST_WB;
	wire REGWRITE_WB, MEMTOREG_WB;	
	wire [15:0] REG3WR_WB;
	wire [1:0] ALU_CNTRL_EX;
	wire [15:0] OPR1, OPR2, OPR_BR_1, OPR_BR_2, RESULT_BR_NPC;
	wire [16:0] RESULT;
	wire [15:0] PC_READ, PC_WRITE;
	wire [15:0] IMM6_RD_SIGN_EXT;
	wire [2:0] REG3ADD_FINAL_RD;
	wire PC_REGREAD_ID, PC_REGREAD_RD, PC_REGREAD_EX, PC_REGREAD_MEM, NPC_CNTRL_MEM;
	wire [3:0] ALUOP_MEM, ALUOP_WB;
	wire [1:0] CZ_MEM, CZ_WB, PREV_CZ_WB;
	wire REGWRITE_WB_FINAL;
	wire [1:0] IRLAST_ID, IRLAST_RD, IRLAST_EX, IRLAST_MEM, IRLAST_WB;
	wire [8:0] IMM9_ID, IMM9_RD, IMM9_EX;
	wire [15:0] IMM9_0_PAD_EX, IMM9_0_PAD_MEM, IMM9_0_PAD_ALURSLT_MEM, IMM9_0_PAD_WB; 
	wire LHI_REG_ID, LHI_REG_RD, LHI_REG_EX;

	
	//IF_stage
	
	instr_mem instrmem_dut(PC_READ,IR_IF);
	assign PC_IF = PC_READ;
	
	ALU_PC alupc_dut(PC_READ,16'h0001,NPC_IF);
	
	IF_ID_reg ifid_reg(clk,IR_IF,NPC_IF,PC_IF,IR_ID,NPC_ID,PC_ID);
	
	assign PC_WRITE = (NPC_CNTRL_MEM != 1'b1) ? NPC_IF : RESULT_BR_NPC;
	
	//ID_stage
	
	controller cntrl (IR_ID,REGWRITE_ID,MEMTOREG_ID,MEMREAD_ID,MEMWRITE_ID,BRANCH_ID,ALUOP_ID,ALUSRC_ID,REGDEST_ID, PC_REGREAD_ID, IRLAST_ID, LHI_REG_ID);
	
	assign REG1ADD_ID = IR_ID[11:9];
	assign REG2ADD_ID = IR_ID[8:6];
	assign IMM6_ID = IR_ID[5:0];
	assign REG3ADD_ID = IR_ID[5:3];
	assign IMM9_ID = IR_ID[8:0];
	
	ID_RD_reg idrd_reg (clk,NPC_ID,REG1ADD_ID, REG2ADD_ID, REG3ADD_ID, IMM6_ID, PC_ID, IMM9_ID,
									NPC_RD, REG1ADD_RD, REG2ADD_RD, REG3ADD_RD, IMM6_RD, PC_RD, IMM9_RD,
									REGWRITE_ID,MEMTOREG_ID,MEMREAD_ID,MEMWRITE_ID,BRANCH_ID,ALUOP_ID,ALUSRC_ID,REGDEST_ID,PC_REGREAD_ID, IRLAST_ID, LHI_REG_ID, 
									REGWRITE_RD,MEMTOREG_RD,MEMREAD_RD,MEMWRITE_RD,BRANCH_RD,ALUOP_RD,ALUSRC_RD,REGDEST_RD,PC_REGREAD_RD, IRLAST_RD, LHI_REG_RD);
	//RD_stage
	
	reg_file regfile(clk, REG1ADD_RD, REG2ADD_RD, REGDST_WB, PC_WRITE, PC_READ, REGWRITE_WB_FINAL, 
								REG3WR_WB, REG1DATA_RD, REG2DATA_RD, PC_REGREAD_RD);
	
	assign IMM6_RD_SIGN_EXT = {10'b0000000000, IMM6_RD};
	assign REG3ADD_FINAL_RD = (REGDEST_RD==1'b1) ? REG2ADD_RD : REG3ADD_RD;
	
	RD_EX_reg rdex_reg (clk,NPC_RD, REG1DATA_RD, REG2DATA_RD, IMM6_RD_SIGN_EXT, REG3ADD_FINAL_RD, PC_RD, IMM9_RD,
									NPC_EX, REG1DATA_EX, REG2DATA_EX, IMM6_EX, REGDST_EX, PC_EX, IMM9_EX,
									REGWRITE_RD,MEMTOREG_RD,MEMREAD_RD,MEMWRITE_RD,BRANCH_RD,ALUOP_RD,ALUSRC_RD,PC_REGREAD_RD, IRLAST_RD, LHI_REG_RD,
									REGWRITE_EX,MEMTOREG_EX,MEMREAD_EX,MEMWRITE_EX,BRANCH_EX,ALUOP_EX,ALUSRC_EX,PC_REGREAD_EX, IRLAST_EX, LHI_REG_EX);
	
	//EX_stage
	
	alu_control alu_cntrl_dut (ALUOP_EX,ALU_CNTRL_EX);
	
	assign OPR2 = ALUSRC_EX[1] ? IMM6_EX : REG2DATA_EX;
	assign OPR1 = ALUSRC_EX[0] ? REG2DATA_EX : REG1DATA_EX;
	
	ALU alu_dut(ALU_CNTRL_EX, OPR1, OPR2, RESULT, ALU_Z_EX);
	
	assign ALU_RESULT_EX = RESULT[15:0];
	assign ALU_C_EX = RESULT[16];
	
	assign OPR_BR_1 = IMM6_EX << 2;
	assign OPR_BR_2 = NPC_EX;
	assign IMM9_0_PAD_EX = {IMM9_EX, 7'b0000000};
	
	ALU_BR alu_br_dut(OPR_BR_1, OPR_BR_2, RESULT_BR_NPC);
	
	EX_MEM_reg exmem_reg(clk,RESULT_BR_NPC, ALU_RESULT_EX, ALU_Z_EX, ALU_C_EX, REG2DATA_EX, REGDST_EX, PC_EX, IMM9_0_PAD_EX,
						NPC_MEM, ALU_RESULT_MEM, ALU_Z_MEM, ALU_C_MEM, REG2DATA_MEM, REGDST_MEM, PC_MEM, IMM9_0_PAD_MEM,
						REGWRITE_EX,MEMTOREG_EX,MEMREAD_EX,MEMWRITE_EX,BRANCH_EX,PC_REGREAD_EX, ALUOP_EX, IRLAST_EX, LHI_REG_EX,
						REGWRITE_MEM,MEMTOREG_MEM,MEMREAD_MEM,MEMWRITE_MEM,BRANCH_MEM,PC_REGREAD_MEM, ALUOP_MEM, IRLAST_MEM, LHI_REG_MEM);
	
	//MEM_stage
	
	data_mem datamem_dut(MEMWRITE_MEM,MEMREAD_MEM,ALU_RESULT_MEM,REG2DATA_MEM,MEMRD_DATA_MEM);
	
	assign NPC_CNTRL_MEM = BRANCH_MEM && ALU_Z_MEM;
	assign CZ_MEM = {ALU_C_MEM, ALU_Z_MEM};
	assign IMM9_0_PAD_ALURSLT_MEM = (LHI_REG_MEM == 1'b1) ? IMM9_0_PAD_MEM : ALU_RESULT_MEM;
		
	MEM_WB_reg memwb_reg(clk, IMM9_0_PAD_ALURSLT_MEM, MEMRD_DATA_MEM, REGDST_MEM, PC_MEM, 
						ALU_RESULT_WB, MEMRD_DATA_WB, REGDST_WB, PC_WB, 
						REGWRITE_MEM,MEMTOREG_MEM, CZ_WB, CZ_MEM, ALUOP_MEM, IRLAST_MEM,
						REGWRITE_WB,MEMTOREG_WB, PREV_CZ_WB, CZ_WB, ALUOP_WB, IRLAST_WB);
	
	//WB_stage
	assign REG3WR_WB = MEMTOREG_WB ? MEMRD_DATA_WB : ALU_RESULT_WB;	
	regwrite_cntrl regwrite_cntrl_dut(IRLAST_WB, PREV_CZ_WB, ALUOP_WB, REGWRITE_WB, REGWRITE_WB_FINAL);
	
endmodule 